library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TB_CLCD IS
END TB_CLCD;

architecture Behavioral  of TB_CLCD is

COMPONENT CLCD
PORT(
	RST : IN STD_LOGIC;
	CLK : IN STD_LOGIC;
	LCD_E : OUT STD_LOGIC;
	LCD_RS : OUT STD_LOGIC;
	LCD_RW : OUT STD_LOGIC;
	LCD_DATA : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	
	);
END COMPONENT;

SIGNAL RST : STD_LOGIC := '1';
SIGNAL CLK : STD_LOGIC := '0';
SIGNAL LCD_E : STD_LOGIC := '0';
SIGNAL LCD_RS : STD_LOGIC := '0';
SIGNAL LCD_RW : STD_LOGIC := '0';
SIGNAL LCD_DATA : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";

BEGIN

PROCESS

BEGIN
	WAIT FOR 10 NS;
	CLK <= NOT CLK;
END PROCESS;

RST <= '1', '0' AFTER 15NS;

U_CLCD : CLCD
PORT MAP (
	RST => RST,
	CLK => CLK,
	LCD_E => LCD_E,
	LCD_RS => LCD_RS,
	LCD_RW => LCD_RW,
	LCD_DATA => LCD_DATA
	);
	
	END Behavioral ;
